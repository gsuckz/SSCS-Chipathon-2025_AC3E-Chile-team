** sch_path: /foss/designs/SSCS-Chipathon-2025_AC3E-Chile-team/xschem/gf180_digital/PD/tb_PD_vto1p1.sch
**.subckt tb_PD_vto1p1
VCC Vdd GND {Vdd}
VSS Vss GND 0
Vg1 VIN_1 VSS PULSE(0 {Vdd} 0 {TR} {TF} {T*D} {T} 0)
C1 V_PWM Vss 10f m=1
Vg3 VIN_2 VSS PULSE(0 {Vdd} {Td} {TR} {TF} {T*D} {T} 0)
x1 Vdd Vss VIN_2 V_PWM VIN_1 PD_vto1p1
Vg2 Vctrl VSS PULSE(0 {Vdd} 0 {TR} {TF} {T*0.615} {T} 0)
**** begin user architecture code


.param Vdd = 5
.param VH = 5
.param Del = 0

.param T = 0.1u
.param TR = 1p
.param TF = 1p
.param DD = 0.615

*Caso 1 - No funciona bien
*.param D = 0.8
*.param Td = 0.03u

*Caso 2 - Funciona bien
*.param D = 0.5
*.param Td = DD*T

*Caso 3 - Funciona bien
*.param D = 0.615
*.param Td = 0.03u

*Caso 4 - No funciona bien
.param D = 0.615
.param Td = 0.08u




.param temp = 27





.save all

.control
set color0 = white
tran 100p 300n
plot v(VIN_1) v(VIN_2)+6 v(V_PWM)+12
plot v(V_PWM) v(Vctrl)+6
.endc

.measure tran tdead_fall
+ TRIG tran1.V(vcn) TD=0u VAL=0.6 FALL=1
+ TARG tran1.V(vcp) TD=0u VAL=0.6 FALL=1

.measure tran t_large_delay
+ TRIG tran1.V(x1.C1) TD=0u VAL=0.6 RISE=1
+ TARG tran1.V(x1.B2) TD=0u VAL=0.6 RISE=1




.include /foss/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/spice/gf180mcu_fd_sc_mcu9t5v0.spice
.include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical

**** end user architecture code
**.ends

* expanding   symbol:  gf180_digital/PD/PD_vto1p1.sym # of pins=5
** sym_path: /foss/designs/SSCS-Chipathon-2025_AC3E-Chile-team/xschem/gf180_digital/PD/PD_vto1p1.sym
** sch_path: /foss/designs/SSCS-Chipathon-2025_AC3E-Chile-team/xschem/gf180_digital/PD/PD_vto1p1.sch
.subckt PD_vto1p1 VCC VSS VINS V_PWM VINR
*.iopin V_PWM
*.iopin VCC
*.iopin VSS
*.iopin VINS
*.iopin VINR
C2 VFE1 VSS 100f m=1
C1 VFE1 VSS 100f m=1
x1 V_N net1 V_PWM VCC VCC VSS VSS gf180mcu_fd_sc_mcu9t5v0__nor2_1
x3 VCC VSS VFE1 VINR net2 SPG_vto1p1
x2 VCC VSS VFE1 VINS net1 SPG_vto1p1
x4 net2 V_PWM V_N VCC VCC VSS VSS gf180mcu_fd_sc_mcu9t5v0__nor2_1
.ends


* expanding   symbol:  gf180_digital/SPG/SPG_vto1p1.sym # of pins=5
** sym_path: /foss/designs/SSCS-Chipathon-2025_AC3E-Chile-team/xschem/gf180_digital/SPG/SPG_vto1p1.sym
** sch_path: /foss/designs/SSCS-Chipathon-2025_AC3E-Chile-team/xschem/gf180_digital/SPG/SPG_vto1p1.sch
.subckt SPG_vto1p1 VDDd VSSd VFE VIN VRE
*.iopin VIN
*.iopin VFE
*.iopin VRE
*.iopin VDDd
*.iopin VSSd
x2 predly net2 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x3 vinn predly VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x4 dly8 net1 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x5 VIN vinn VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_2
x6 predly V_gatein VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_8
x1 dly7 dly8 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_8
x8 net2 dly8 VFE VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__and2_1
x7 net1 predly VRE VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__and2_1
x10 VDDd VSSd V_gatein dly7 large_delay_vto1p1
.ends


* expanding   symbol:  gf180_digital/large_delay/large_delay_vto1p1.sym # of pins=4
** sym_path: /foss/designs/SSCS-Chipathon-2025_AC3E-Chile-team/xschem/gf180_digital/large_delay/large_delay_vto1p1.sym
** sch_path: /foss/designs/SSCS-Chipathon-2025_AC3E-Chile-team/xschem/gf180_digital/large_delay/large_delay_vto1p1.sch
.subckt large_delay_vto1p1 VDDd VSSd VIN VOUT
*.iopin VIN
*.iopin VOUT
*.iopin VDDd
*.iopin VSSd
x1 VIN VOUT VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__dlya_1
.ends

.GLOBAL GND
.end
